library verilog;
use verilog.vl_types.all;
entity ALU2_vlg_vec_tst is
end ALU2_vlg_vec_tst;
